`timescale 1ns/1ps
module 189_OoO 

 
   






endmodule