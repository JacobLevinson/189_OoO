`timescale 1ns/100ps

module complete_rob import typedefs::*;(
    input logic clk,
    input logic reset,
    input completeStruct complete1,
    input completeStruct complete2,
    input completeStruct complete3,
    input robDispatchStruct dispatch,
    output forwardStruct forwarding,
    output 
);



endmodule