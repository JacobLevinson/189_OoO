module rename (
    input logic clk,
    
);



endmodule

